module main

fn reverse_string(str string) string {
    return str.reverse()
}